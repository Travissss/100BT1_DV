//////////////////////////////////////////////////////////////////////////////////
// Engineer: 		Travis
// 
// Create Date: 	02/17/2021 Wed 19:46
// Filename: 		chnl_pkg.sv
// class Name: 		chnl_pkg
// Project Name: 	mcdf
// Revision 0.01 - File Created 
// Additional Comments:
// -------------------------------------------------------------------------------
// 	-> VIP for mcdf channel
//////////////////////////////////////////////////////////////////////////////////

`ifndef MCDF_CHNL_SV
`define MCDF_CHNL_SV

package chnl_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"



	
endpackage

`endif